library verilog;
use verilog.vl_types.all;
entity test_ulaControl is
end test_ulaControl;
