library verilog;
use verilog.vl_types.all;
entity test_memoria is
end test_memoria;
