library verilog;
use verilog.vl_types.all;
entity test_registradores is
end test_registradores;
