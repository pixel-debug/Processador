library verilog;
use verilog.vl_types.all;
entity test_ula is
end test_ula;
