library verilog;
use verilog.vl_types.all;
entity test_dados is
end test_dados;
