library verilog;
use verilog.vl_types.all;
entity test_memoria_dados is
end test_memoria_dados;
