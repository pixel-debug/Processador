library verilog;
use verilog.vl_types.all;
entity test_controle is
end test_controle;
