library verilog;
use verilog.vl_types.all;
entity test_adder is
end test_adder;
