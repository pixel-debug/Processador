library verilog;
use verilog.vl_types.all;
entity test_jumper is
end test_jumper;
