library verilog;
use verilog.vl_types.all;
entity test_processador is
end test_processador;
