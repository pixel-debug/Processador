library verilog;
use verilog.vl_types.all;
entity test_extensor is
end test_extensor;
