library verilog;
use verilog.vl_types.all;
entity test_pc is
end test_pc;
